
-----------------------------------------
-- Definition of Hybrid Carry Look Ahead(CLA)
-- and Ripple Carry Adder(RCA) 4 Bits
-----------------------------------------

Library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.MTNCL_gates.all;
use work.ncl_signals.all;
use ieee.math_real.all;

entity SYNC_SF_Core_wo_input is
generic(bitwidth: in integer := 8);
	port(
		clk  				: in std_logic;
		reset  				: in std_logic;
		parallelism_en  	: in std_logic;
		id  				: in std_logic;
		pixel_out   			: out std_logic_vector(2*bitwidth-1 downto 0)
	);
end;

architecture arch of SYNC_SF_Core_wo_input is

component SYNC_Weighted_Box_Filter_W_reg is
    generic(bitwidth: in integer := 8);
    port(
    		clk : in std_logic;
			input    	: in  std_logic_vector(bitwidth-1 downto 0);
			reset  		: in std_logic;
			output   	: out std_logic_vector((bitwidth-1) downto 0)
      );
  end component;

component SYNC_SF_Data_Loader_wo_input is
    generic(bitwidth: in integer := 8);
    port(
    		clk : in std_logic;
			inputMUX    	: in  std_logic_vector(4096*bitwidth-1 downto 0);
			reset  		: in std_logic;
			parallelism_en : in std_logic;
			id: in std_logic;
			clk_out : out std_logic;
			output   	: out std_logic_vector((2*bitwidth-1) downto 0)
      );
 end component;

signal clk_out : std_logic;
signal pixels : std_logic_vector (2*bitwidth-1 downto 0);
signal pixel_in : std_logic_vector (4096*bitwidth-1 downto 0);

begin

pixel_in <= "10100000100111101001110010011010100111101010101010100111100000100101111101100111011010110110110001101100011100100111101101111111100000111000010010000010100000111000011010000110100001101000010110000111100001101000010110000011100001001000010010000101100001011000010010000010100000011000000110000001011111110111101001101101011110011001011010011110100110001001101110011011100110011001100110011100100110111011000111011100101110110110110001110101011110100111101001111010011111000111101101111101011111010111110110000101100111011001110110011011100110101010001010101010101000100111111001011100011001000110101001101001011010000111000001111001011111101000000110000011100000101000001010000011100001011000010010000100100001001000010010000100100000101000001110000011100001001000001110000011100000101000000010000000100000001000000001111010011100010110111110001011100111011001110110011101100111101001101110011010100110101001100110011100110010111101100010001101011011000111100001111001011110010111101101111100011111101000001101100001001100101001101110011101100111001001110110100110101001101001111010000000010111010110010001101010011001110110011101110001011110000111111010000010100000111000001010000010100000111000010010000100100001011000010010000100100000111000001110000010100000101000011010000101100000111000001010000001011111111000000010000000011111010111010101101011011111101001101010100010101000011010000110011110100110111001100110011001100101001010101111011011110001000111000101110010011110100111101001111100100000011000011001011110001100000011000010011101100111111001111010100100101001101010000010011111011111110101101001100100011010110110100001101000011100000111100101111101100000011000000110000000100000101000001110000011100000011000001110000101011111110111110001111111011111110111111110000001100000101000010010000001100000000111111001111111100000000111110101110101011011000111101110010110101000001010000010011110100111101001110010011010100110101001011010010101110001001101111110011111011011000111100101111010011111001000010101011100001011110010111000110101100111111010000110100100101001111010010010011111100111110111110101011001011001000110100101100111011010000111000101111000011110110111111110000000011111101000000010000001100000011000001010000010100000100111111001111001011110100111100101111000011111101000001010000010100000001000000001111110011111110111111101111100011101010110111001111001100100001001101110011110100111011001110110011100100111001001101110011001100100001010000111011010110101000111110101101111011110111000001001011001001011000011010000110100001100111010000110100011101001011001110110011110101000001001111101111101010110000110010001101001011001110110100001110001011110000111101101111110011111010111111010000000100000001000000110000001100000001000000010000010100000101000011110001100100010001000000101111011011111000111111110000001011111110111111101111111011111000111010001101111011101111000110010010101100110101001101110011010100110101001101010011001100101011001000010001111110000001110001110110000011010110111100001011010001011000011001100111010001100110010111110100001101001111001101110001100100111011010010010100000011111100101011101100001011010000110100001101001011100100111100101111100011111100111111110000001100000001000000010000001100000011000001110001111100100011001101010100111101100101011000110110000101001101000110101111000011111011000000001111111011111010111100101110100011011100111011110001101100100011001011010011010100110011001100010010111100100111000111110001110100011001001101111010101110111101001001101010100001010100010111100110111001101100011000000101111101001001010011010000100011111101010000110100110101000110111111101010010010111010110001101100101011010010111000001110111011110010111110001111110011111100111111110000101100010010111111110000101100010101001000110011000101000011010101010110001101101111011111011000010101010010111111101110101011110110111101101110101011100000110101001110101100011101001001010010011100101101001011110010010100100001001000110001110100011001000110110001010101100101110101010101101001010100010111000110110001100110011001000110000001100011010110010011000011000100111011110100010101001101010000101111100010011110101101001100010011001000110011101101101011100100111010101111010011111000111110010000000011110000111101001111011100000011000001110001000100011111001101110101010101100101011100010111100110000001100100010111010100010010110100001110001011100110110111001101000011101001001000010010101100100101000111110010010100100011000111110010001100011111000111010001111100011111001101110111110010101100010100000110100001101010011001000110001001100110010101110100110011110110101000101111001101000111010100010011111011110110100111101011100011001000110010001100110011011010111001101110101011101110111101010000001011110010110111101110101011111011000000010000101100001111000101010010101101001001011001110111010101111101100000111000001110001011100101010101001011010110110100101101001011001100111001010010011100111001001010101111110011111111001010010010001100100011000111110001111100100101001011010010111010011110010011100110011001101000011000100110100001101100011010101011010100100010101111001010101011110111010001010101000100111110111101001010000010110110110001101100101011001100110110101110010011101100111100101111100011110100110111001110011011110000111100001111100100001001000011110001001100100011010001110110110101110001011011010111111110010101101000011010010111000011010100001011001011000100110001001110001100100101001110010011001011101000101010110000110100101001001000110001111100100001001000110011011011001000010011000110010001101100011000100110010001100110100000101011000100101010110111101010111010110000111101010100000101010001001111101111001010100010101110101100011011001000110011001101101011101000111011101111001011110100110111101110001011101100111010001110110011111111000100110001101100011011001000010100001101010101011000011000011110011101100110111001010110011011101001111011110100010000100111101011011011011111001001110011011100110010111100000110111011001111001001010010010100011111001000010011000100000000011001000101111001101110011001000110100001100010011101101011101100011011001010101011001010111000101100101111000100111101010011010100000011110010101000101011101011000110110001101100101011010110111010001110110011111000111010001101111011100010111010001110111011111111000010110001010100011011000100110001011100110011010110111000011110010011100011111000110110010011100110011001111110101001101011010001111010010100110101110010010100110111001101001111010001100110100000110000000100100111000110010010010100101010100010000101001001110000011010000110010001100100011001001001101100010001001011010100001010110100101110001011001011110001001111010100101101000000111101101010001010110100110001001100100011001100110110101110011011101011000100001101010011011110111000101110100011110111000011010001010100010101000100101111101100011001011000011000001101111111011110111000011110010111100110011001101110011011100111011010101110111000111001001011110100100011001101110011011011110110011100000100111010011101000111010010111100101100110001100101010001101000011011100110100001101000011001000111010100000001001000110011101101000110101101101011011010101100111011010011110101001001010000001111100010011110101100001100001011000100110011001101100011011010111111010010001011001100110111101110001011101111000001010000110100001101000010101111010100011111011001110110111101101111011100011000001110001001100011011000111110010011100101011001101110011111101101010111100010111001000111010011010100110110111110000110111001000100110010011000001110100101100010000111110001011100011011100110111001101010011010100110001011011101001010010011010101000001001111001011011010111100101101101110110100111101010100010100000011110010100101101010111011000100110001101100110011010110110110010010101100011010110010101101110011100100111110001111101011111111000000001111001100110001010111010101100101011111011001110111100101111011011110111000000110001001100100011001001110010101100110011001110110101111000101010000111100111011001101101110001001100100111101011000011110101001101100011100010010111110010110000110110001100010011000100110010010101101001010010011000101000001001111010011100011000100110001101100000011101101001111010101001101000110111110001010000010110100110010101100110011001110110111001101101101000111000001001100011011010110111010101111010011111000111111101111010100101001010001010100011101011011011010010110110101101101011000110110111110000001100010011000101110000111011111011001000110010101100110111001010100111101001011110010010011111011010000011001010110011111100111011001101110111110110010000101101001101000010111100110001001101101000011110011001101000001001110110011100100111000110010101100101011000100111101010011110101010101010100001111111010100100101110001100101011001100110010101101011011011001010101001111111011001100110100001101110011110000111101001111011100011111001011010010100101000101010110010101110101011111010101110110000101101001011011010111011101111101011011110111011110000111100001111000011110001011011101110011011101011101100001111001100110011011100101111001011110100111101100001010000001100000011000100110000001100110110011110011000100111001001111110011101100110111001101001100100011000110110001001111010101000011010111010101010100000000101000001011011011001000110010001100011011001110110111110110111100010010110110101101010011100000111100001111011100011111001000010001011100101101001110110100111101010011010100010101101101011101010110110110010101101101011001110111001101111101011101010110110101101111011001010111011101111111100100111001010110010011100100011001100110001001101010011000110001110000011000100110001001011110100111010010001100110011010000010011111100111011001101110011100011000100110000101100000011110011010001010101101101010011000000001010001010111000110001101100011011000110110010101110010101110001001100001111110011010000110110001110110100010101000101110000110100101001001001110010101100111101010011010101010101010101010101110100110101001111010110010110001101101111011001110110000101010011010110010110111110000011100011111000111110001101100011111001100110000111010011110111110100100010010101100110010001011110011100001110111100110001001111110100000100111111001111010011101100111000110000001011111011000000111110010100010101011001010100010000010010100100101110101100011011000100110010001100001011100101011100110011110100010100110110001101111100001111000011010000010100011111000110110010000100101011001101110100001101000101001111010100001101000011010010110101000101010101010101010100101101001001010110110111010110000111100001111000010110000111100100111001010110011101010111110011010101011100101101000101011001100110010111101011010100101101001101010100000100111011001111010011101100111011001110001100010011000010110010001111110101000111010110110101010100000110101000101011011011000100110001001100011010111100111001111000011101010001001011101111010011111001000001001111111100010101000011110000110100011101001001010001000011111111000000010001101100010011001011110011010100110011000100010001110101000011011000110111111110000111011111111000001110001101100100111001100110101001011110110000000011111111010100100110010001011110011010000111010011111111001100010011110100111011001110010011100100111001001101110011010011001000110001101100111100000011010010010101110101010111000010001001111010110100110001001100100011001000101111101101101110010001011001010001100011111010111011001111000100010001000001110000001100001101000101110000101011111000110100101011001100001010110110001011100010110100100000000111001011111111011010111000001110000111100001011000001110001101100101011001111101111101001100101101010011001101010101001101001001010100011000100101110010100011001001110011100101000001001111010011100100110111001101010011010100110010110100001100101011010001000000110100011101011011010101010000100010100000101101001100010011000110110001101100001011000001011111010111001100001101000001101110001100001001000001001111111100000111000100010000000011101110110010101010000010001100110001001010101010101100011111000110100011101111010101110111101110000011011111010111111110000011100101011000000101000010110101101100010100000101010111101100111001011010011001000110011001101100111011010011001101000111010000110100000100111101001110010011011100110101001100001101011011001110110010101111110101000011010110010101010100001100101000001011010011000010110001101100011011001000101101110100000110001011001110101111101011111100111111001111011011111101000000001111100011010100100111101000001001100100100111001001100010101110100010001001100100000111011001010111001101101101011010110110111101111101100000010010101011011000111011010010101101010001011011101101000001010100011011000110001001100010100101010001111100111011010010110100100101000011001111010011100100110111001101010011001011011000110011101100011011110111010001110101101101010111000011001001110010110000110000001100010011000100110011001100101011101101100010010101101011111110111110101111011011111010111111101111001010110000100111000111101010001000011100001000011001111010100110001011000011110011011001111000001101101011011001010101111101101111011111110101100010101100110010001111010100111101010101001011011001010010011010000110110001011110011001101100101100100001010010110100011101000111010001010011111100111101001110110011011100110010110110001101000011000000111010110100001101011011010110110000111010011100101011001100000011000100110001101100111011011100110000110101111101111100111111001110100011111000111111101111000010110010100010001010000001110010100101000111111001100110011011001001000011010101001110010111001101100011010111110101101101100011011111011000011110000110111101001001110011011011001010001001111001001010011010100111010001100110010111001000001011110101001001010101000101001011010010010100010101000011010000010011110100111001001100001101010011010000101111101110011101000001010111010101100100010000100111101010111011000100110010001100011011010010111000101100111101010111010101101101110011101010111101101111011010100010011111000101111010000110100011001000100010101000010101000111011011101011001000110110011101101101010010110101010101010011011101111000111110010011100111010010110001110010101000010001100001111000010111000111001001111000011000000101101010110111000101010010111100111111010001110100010101000101010001010100000100111101001110110010111011010010110011101011111011100111010000010101110101011011000101001010010010110010110011001100111011001000110111001110111011011111000111110011000011011100111111001110010010010010011100100111100001101010011010100111110010100000100111000110101100000001010101110100001101100011011000010100010101000011011001011000011110010001100111011010101101100010100011000110100100001100100010000110100001111000011101000101111001101000111011110010101100111011001011010010111100110011001101110011111100111111001110110011010100101110110100001100100010111010111001010100000101011111010110110001001010100110101101101100101011001110110011101101110011101010111010001111010100001110111111001111111010011100011110100110011010000010011101100110110001110110100000001000000011101011001111110110101101010111010111110100101101000101010101110110100110000101100011111001100110101011100011001100001001010110111100101001110001101100011111000110111001100000100101010001010100111101010001010011111100111101001101010010011100100111001001110010110100110001001100001100110011001000101111101110001101000001011000010101110100010010101001001011001011001100110011001100111011011100111010110000001011100000110011110000111011000010100000101000110001101100100001000110011001110000100001100111001010110011001110110101000101101001011001110000110100001011001011110110000101100011011101111000001110001111101001011000000010111110010011101101011010111100011101100111111001101000011000101100110100100001010000110011111101000001010001110100001100110101001010110010001100100001000111110001111011001100110011101011110011100001010000010110000101100001000101101010100010110110110011001100110011001010110100101111000100100110110110101011100011001100100100101001000010011010011100000111011001101110011001000111110010001111001010110111000101100111010011110000010011110100110110101011101011111101010011010110100110000001011110110010001011010100101011000101110010111110110100100111100001110100011001100111011011110101001010110100001100111011001110010011100100111101001101010011010100110111001011010010000100001110110001101100010010110000110101110100001101100011011000010001100010100010101100101100100011000110101111110000000100101011001100110000001010010010100011001010011010110000011110001000001001100110100011100110100001011000111110110110010110001101001101101001010001110100011111001010000010100000111110010010000101100001100011001111000010001110100000100111100001011110101100001110010001111010011010100110000010001111000101010011011100111011001101010011010100110101001101110011001100110011001100110010100100011111000011101100010010111110101000101100101101000001011001010110000100010110101010001011101011001000110010001010010100000001010111101111110010000010011111101000100010010010110001100110010001101110011101100101111001011100101001010011111101111111011001001101001010000000100110001100000101101110110110101110010100001111011100110101011010010000110011101101111001011010010110101010111011110000100001100110011001011110110000110010100100111011001101010010111100110001001100110011001100101111001010010010001100010011000010110001111011001100110000101010001011001001010000110110100101101001000110101011001011000110110111101011100011001101000101110000100010001010101001001000101010001000101100101110010010001010010110000110010001011000011001110000110101110011010110101111110100010001000000101110101100010111010100110010101011110111000001110111110101011101000000010000110010111100011101000110001010101101000000001000010001100000011100101111001100101101001101110011001100101111001100110011000100110001001001010001100100010001001001010101000101101110110010001011010010010100101110110100000101101001011010110010000010110000110001001101101011111101000010101011011001101110100010001101011010001010100001001011101011100010100110100101100001100000010101101100001101011001011000001101101100000101001100010011110100110001001011010011110100110101000011010000001101101011100011110011011100000000110110001001101001100010101000010001000001111010010111001000100100001111001101010011010100101111001011110010110100101101001001110001101100010001010010010111101101111111011110101011011010100110100010001011001100111101011001110110100100011110101011101100001011110011000001001101011010011000100010001100111010111100011000000111010010110110101101001100001001101110010101101000010100011111011100001011110011010111000010110010111101010001011000010110000101011011001110010001101100000001010101111001110101001001000110110000000010101000011011001001000100010100011100000101100010110011001000010011101100110011001011110010111100101001001001010001110100001111010010111000100110000111011111011000001010011110100110001000000010110001001111010110001101100011000111101010111011000100111001101101101010111000101001001001011011001010100100000110010001100010011101000110100011100100101000000100100011001011011100001110101001111000111011010000101100100101010001010110000101100011010100110011000100011011000000010100100110011101010001010010000100000010100110000110110010000011000101100111110001100010110111110011011100111011001100010010110100100111001001010010001100001111001011011000001110000011100001111000111110010100100111001001010001110110101010010011100101011101010111110001111010101000110110001111111010111110110010101010010010100110110111101010001001100110010101101000110010100011000000001010101001101001001000110100001001011110100010101110001100001001000111110011011101001011010100010100100100100001000001101111100100110011100111110100010100100000111110000111101001111000011101110001001010010010011011110000011100111101001110010011000100101101001001110010001100011001000100110110100110000101100001011001100110100001100101101010010010010110011011001001110100111001011000010110001100011110101011101101011011101000101010101011110010100000101010101101100010101000011001000101101010011100110100001001101001011100110111110100000010011000010101101001111011011101000001010001011100101011001101010100000100111101000010110000001100000001001000011001100101000001000111001101011001011110100000000110101100000100101011001000110100100111001110110011000100101101001011010010100100100011000100010011100110000111100001011001011110011111100111011001110010100100100110100111110010111011001111110101111101100011001001001011100011000100110101001010100010110010101001001010000011001110110110000111001001111010011011001010001001011010101000110110011011100100010100000110110010110010111000010000001100010101001001110011000100111011001110110001010011110000110110110000000101100101001100110001001010011000010111001000011001100100111010001100101011000011001101010011010100101101001011010010101100100101000111110000111101011111100010111000111110011011100111111010000110011100100111001001100010001010111000110100001101011001011001010010100010101100101110101110001010010000101000001001100010011010110010101111000010011000101110000110110010100110111111101111101100001000011010000110101001110100110001101110100100000001000100010001111100101001001101010011101100101111000110010010111101010111011001010010101011110000011010000110110010010100011011001100010011100100111101110011011100110101001011010010101100100111001000110001101100010111011101011000111110011101100111011010000110100011101001001001001010001110100001001110010101000011010101110110011100101010101010001100100011100100101001001010011001111010100011001010001011000100111010001001000010010011000111010011001011100000100010000110001001110110011100001100000011100111000000110001000100011001000110010010100100101111001011010011001101110101100010110110010100011110101011000101101001110110100110000110111010100100111111110001010100110101001100110010101100101011001001010010001100010111001000011000000110011011100111111001111110100001101001011010011001111100100000101000011011100011010001110101111101101001001010001011100011010110110110001000110010001000011111101011001010110010101001101100111010110101001110010101101011101110101000100110010001101000011111000111001010101000110101010000001100001001000110010001101011110100111101010000010100000001000101010010000100001100111111000110111001100010011111101001100001110100100011110001000100100101001101110011000100101001001010010010010100100011000100010010010110001101101000111001111110100011101001111010101110101000011100100111110010001010111010110100100101100011011010010010111011010010110100101101101010001100011011101000111011010100101111101100000010110010111111110100010100100100111000000110100001100010011010000111101001111000100101001011110011110010111110110000111100100011000010001110110011110101000101110011011100100111000110001010110001011010011000100111110010011000100000101000100100100011001011110011011100110011001011010010101100100101001000110000110100110001101000011010100110100101101001111010101110100111101000100110110001101100100011001110001100111111011001010110100100101100101010001110000010101110101000000111010010011000111100101100110010111110111001010000001101000001000111100111110001101100011010100110110001111010011110001000101010011100110101001110110100000001000101010001101100001011000000010000101100011001001010001111010001100100011000100110101001111010101000001000100010001011001010110011001100110101001100110011001100101101001001110001111100000101001101011010111110101011101010111010101110100011100111111001110001100110011000101010011011101001001101110110001101100111001010001010100011001100101000101000100001110100100001101110001011101110110110101101010011011001001101001010000001011110011100000110100001101010011011100111010001110100100000001001111011010000111110110001000100011001001000110010111101000001001111010010011010010110010110100110111001110000100000001010100010010000100010110010101100110111001110010011001100101111001011110010011100011100111110110011100110110111101011011010101110101001101001011010011110101000011000000110000010100000111011010011101101100001011001010010101010100010101100001000110010001100011101100111100011001000101010001111000011110110111101101011011001100110011010100111011001101100011010100110010001110000011101000111111001110110100000101100011011110111000100110010110101001001010100110100100011111110011010000110101001111000011011001000111010110000100110001001010100101101001011010011000100101111001011010010101100100011000101001111011101010101101110111010100110101011101010011010000110000101001101100110001001010100100000101101110100111101010111010110000100100010111001001100100001111110100010100111100001100100111010101011001010111010111011110000110011100110100101000110001010000100011011100110101001100110011010000111100001110110100010001001111011001000111010110000001100100001001101110100000101000001001000101010011001101110011010100110100010010010101101001010001010100101001000101111001011111001000001110001010100100001000111010000111011110111011110111011000110100101101001011001100100101100100101000110011010100110011100000111000010101011001011110101100101011101001111101101011010100110011001001000010001111010100010101011010011011010110100101101011011010100111000001111101010000010011111100111001001101010011001100110011001110000011100101000010011011111000001010000100100010001000111110010001100100101010100111000100110001001001110001011001001010010100011001010111010011100101011010001101100000000111101001110011011011010110111101110100011101010111001111000001110100001101000011001110100100100011111000111000010100001000100001101100010001110100001010010000101010111010111010010111011110000100010100100111010011100100110001010111010000100101111101100010010110000111010010000001011001010101101100111011001110100011011100110101001110000011100001000000001111110110101101111100100000001000101010001100100010111001011110101110101111101100010011001111110011011000001000111110010011000100011101010110100100101001000110001101100001100111101101101111011000110110111001100110101111001101010011010001100100010100001101001001010101110101011110000010100101100110101101000010100100011011000010101110101000111000000100110001001100010100000101000111010000110100000101001010010001110100111001110000100001110110100101101111010001000011100000111010001101110011101100111011010100110100001101101010011110111000010110001100100011001001000010011110101010001011001110111001110000111100111111011010100100010011100101000000010110011001010010010100100100011000111010001001100000100111100101111011100000111100110111011000101110110101000001010000010111110110011001011101010010111001110110001100010001001001000110110010101100001010000001101001001010010011011000110110001101110100110100110010010000010100110001010010010111110111110001111110011000100110000000110010001110100011001100111011001101100110010001001000011001011000001010000111100011011000110110010010100110111010001110101100101101011011111111001001110100111101110001101010001010110101111010010011100100101001000110001110100010111000011001111111100001001010011111010110110101101001000001010010011000100110101101100001011001010010111010010101100101100011111110001111101101001011001010011101011001010010111000110110001011100100010001010000001100100011110001000010010111010101100001110111011110110101011101101010001100110011111100110100001101100011101101101001010011000110100010000100100010001000101110001100100100101001011110011111101010001011000110111100110001111100111111011101101110010010101001100010100101101001001110010001100011001000100010000010100000001010110111001100110110011100010101101101010111000110110101100011011000000110011100100110100010111001100100111111100011101011001110110011100111110101100100110001001011100010111001010111010001100011011000110010001100110100101101011011011101101000001010000000011000100011100100111100001101110011010001010000011110010101001101101100100001111000101010001001100010111000111110010101100111001010010010101110101110101100011011001110110101011101101101001111011001101001100010010010100011101000101110000110011111001001001111010101110101011101101010100011010111100110010001101110010111110110011101100000001000111000010010011111010001011000101110110010101100001001111001011010001011100010111100110111010000110100000100110111001100000011100000111110010100101000000101101001010111110101010001010011010011100011100000111000011001110111111001010011011101001000011110001101100010101000100010001100100100101001101010100000101010011011011111000010110011001101000111011110100000100110111010010111100011111000110010001011100001100111101110100001110101011101010111001011100001000110010001101000011001000110001001100100010110000010001101110101101000010100110110001000101100101011001010100001010111110010110000110101001110010011011100111011001101100011010000111010010001110101010001110011011001110101011100110110001111000100000100110100010001110111010001111000010101011000000110001100100011011000101110001000100010101001000110011000100111101010010110110001110000001100100111001111110110011011001101111111100100011001000110010001100011011000100010000011100101011011110011010110101101100111001001100011010111100101101101100101010111100101111000100010011010101010001101010111100001011011000110110011101000000110011100110010001101100011001000111010001111100011100100110010001110110100111001010000010010110100111101110010001110110011000100101110001100110101101101111011011000110101111110001001100011011000111110001101100010101000100110001111100101101001101010100000101010111011101011000101110011111101010111010011100000010101111001110001100000101000101010001101100100111000100110100000110110001010000101100010010111000101010101100010010111110110000001010000001000000110001010101101011000101000000010101111101100111001110101100010001101010010110100110111001110010011110000111001001011110011010101001101011101000101001001010001010000000011000100101101001010110100011001110000011100100100100101111000100010011000110010001110100011101000101110001000100011001001001010010111100111111010011110110100110000101100110111010011110111001000010101010000010100110100111101001111010111011000101010011010101101111100111101110011010010110101010001011101010111110110000001100000001111010100010101101100101100110111001001111111101011111011010010011010010111100011000100110011001101010011010000111011001111000011000100110011001101010101101001111100011000000011000100101101001010000011001101100000011101100100101101011100100010001000101010001011100011101001000010001101100010011000101110001101100101001001101010100010101011111011110111001001110100001101101010101010011000000110011001010110001111100010011001111000101111111100101010011011010000100100011101011010011000000101010101100111010110000011101101011011011111111011000001111110011111111010111010110111100110000101100100110000001100110011010000110010001111000100001100111001001110110100000001000011011001100101010000101111001010100010101101001011010111110100101101010011011111101000011110001011100010111000110110010000100011111000110110001100100011001001000010010110100111111010100010110101110000111100111011010111110001110110010101101001011001000101011001000010100000011100110010010100010010000011111001010100011000100100110101011100011011000101000001000010010000110110111010101000100001010111111110101111101110001001101001000101001011110011011100111011001110000100000001001000010101010011111101000100010010110110101101001111001011000010110000110001010001000101000001100111011111001000000110000100100010011000101010001101100100001001001010010001100011101000110110001111100101011001110010100101101100011011110011001001110101001101011001110110010111100110100101100110011010000111110010001001010100100100100101010001011001000100111001001100011011110110011101000101001110100011011001010101101100111001111010000010101011111011100110010000001110110011000100111000001111100011110001000011001111110110001001001010010001110100011101010111010100100010110000110000010010110110100101110110011111010111111110000001100000111000011110001001100011001000111010010010100100101001001010010001100100101001010110011010101000101010110010110111110000111100111111011000100011110101010001101100011101000111011001110000011001010110100101011011010111010101000101001001011001100111010101010011001110100011100000110000010010101011110110110010100001011010111010111000100010010011011100110010001111000100010001000100010100110100010001010101010101100100111100111110010000010101010001000111010001110110001101110100011110100111111001111111100000111000010010000111100001111000101010001110100100101001000110010011100101101001010110010111100111001010001010101000101100111011111111001000110101001011000101011000011000100111010001111110011110011000000101110000010110000101010101010011011000000111111001011110001101110011100101011000";

sf_data_loader_instance : SYNC_SF_Data_Loader_wo_input
 generic map(bitwidth => bitwidth)
  port map(
  					clk => clk,
				    inputMUX => pixel_in,
				    reset => reset,
				    parallelism_en => parallelism_en,
				    id => id,
				    clk_out => clk_out,
				    output => pixels
    );

box_filter_instance_a: SYNC_Weighted_Box_Filter_W_reg
 generic map(bitwidth => bitwidth)
  port map(
  					clk => clk_out,
				    input => pixels(bitwidth-1 downto 0),
				    reset => reset,
				    output => pixel_out (bitwidth-1 downto 0)
    );   

box_filter_instance_b: SYNC_Weighted_Box_Filter_W_reg
 generic map(bitwidth => bitwidth)
  port map(
  					clk => clk_out,
				    input => pixels(2*bitwidth-1 downto bitwidth),
				    reset => reset,
				    output => pixel_out (2*bitwidth-1 downto bitwidth)
    );  

end arch;
